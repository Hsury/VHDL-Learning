--流程控制模块 2017/04/27
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FLOW_CTRL IS
	PORT (CLK_50MHZ : IN STD_LOGIC;	--50MHz时钟
	      KEY_MASTER : IN STD_LOGIC;	--主持人按键
	      KEY_CLIENT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);	--客户端按键
	      LED : OUT STD_LOGIC_VECTOR (3 DOWNTO 0));	--状态指示灯
END FLOW_CTRL;

ARCHITECTURE BEHAV OF FLOW_CTRL IS
	TYPE STATES IS (S0, S1);
	SIGNAL ST : STATES;
	SIGNAL LOCK : STD_LOGIC;
BEGIN
	PROCESS (CLK_50MHZ) --Mealy型有限状态机的状态切换及控制进程
	BEGIN
		IF RISING_EDGE (CLK_50MHZ) THEN
			CASE ST IS
				WHEN S0 => IF KEY_MASTER /= '1' THEN	ST <= S1;	END IF;
				WHEN S1 => IF KEY_CLIENT /= "111" THEN	ST <= S0;	END IF;
				WHEN OTHERS => ST <= S0;
			END CASE;
		END IF;
	END PROCESS;
	
	PROCESS (ST)	--Mealy型有限状态机的输出控制进程
	BEGIN
		CASE ST IS
			WHEN S0 => LOCK <= '1';	LED(3) <= '0';
			WHEN S1 => LOCK <= '0';	LED(3) <= '1';
			WHEN OTHERS => LOCK <= '1';	LED(3) <= '0';
		END CASE;
	END PROCESS;
	
	PROCESS (LOCK, KEY_CLIENT)	--注意: 锁存器(Latch, 电平触发型寄存器)需将输入信号加入信号敏感列表!
	BEGIN
		IF LOCK = '0' THEN
			LED(2 DOWNTO 0) <= NOT KEY_CLIENT;
		END IF;
	END PROCESS;
END BEHAV;