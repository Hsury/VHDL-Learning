--按键消抖模块 2017/04/11
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY KEY_SCAN IS
	GENERIC (KEY_TRIGGER : STD_LOGIC := '0');	--配置按键触发电平
	PORT (CLK_1KHZ : IN STD_LOGIC;	--1KHz时钟
	      KEY_IN : IN STD_LOGIC;	--按键输入
	      KEY_OUT : OUT STD_LOGIC := NOT KEY_TRIGGER);	--按键输出
END KEY_SCAN;

ARCHITECTURE BEHAV OF KEY_SCAN IS
	SIGNAL CNT_KEY_DOWN, CNT_KEY_UP : INTEGER RANGE 0 TO 9;
BEGIN
	PROCESS (KEY_IN, CLK_1KHZ)
	BEGIN
		IF RISING_EDGE (CLK_1KHZ) THEN
			IF KEY_IN = KEY_TRIGGER THEN
				CNT_KEY_UP <= 0;
				IF CNT_KEY_DOWN < 9 THEN
					CNT_KEY_DOWN <= CNT_KEY_DOWN + 1;
				ELSE
					KEY_OUT <= KEY_TRIGGER;
				END IF;
			ELSE
				CNT_KEY_DOWN <= 0;
				IF CNT_KEY_UP < 9 THEN
					CNT_KEY_UP <= CNT_KEY_UP + 1;
				ELSE
					KEY_OUT <= NOT KEY_TRIGGER;
				END IF;
			END IF;
		END IF;
	END PROCESS;
END BEHAV;