--3-8译码器模块 2017/04/11
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DECODER_3TO8 IS
	PORT (DATA_IN : IN STD_LOGIC_VECTOR (2 DOWNTO 0);	--二进制光标
	      DATA_OUT : OUT BIT_VECTOR (5 DOWNTO 0));	--数码管位
END DECODER_3TO8;

ARCHITECTURE BEHAV OF DECODER_3TO8 IS
BEGIN
	DATA_OUT <= "011111" ROR CONV_INTEGER (DATA_IN);
END BEHAV;