--时钟分频模块 2017/04/27
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FREQ_DIV IS
	PORT (CLK_50MHZ : IN STD_LOGIC;	--50MHz时钟
	      CLK_1KHZ : BUFFER STD_LOGIC);	--1KHz时钟
END FREQ_DIV;

ARCHITECTURE BEHAV OF FREQ_DIV IS
	SIGNAL CNT_1KHZ : INTEGER RANGE 0 TO 5E4 - 1;	--1KHz时钟计数器
BEGIN
	PROCESS (CLK_50MHZ)	--1KHz分频器
	BEGIN
		IF RISING_EDGE (CLK_50MHZ) THEN
			IF CNT_1KHZ = 0 THEN
				CLK_1KHZ <= '1';
				CNT_1KHZ <= CNT_1KHZ + 1;
			ELSIF CNT_1KHZ = 5E4 / 2 THEN
				CLK_1KHZ <= '0';
				CNT_1KHZ <= CNT_1KHZ + 1;
			ELSIF CNT_1KHZ = 5E4 - 1 THEN
				CNT_1KHZ <= 0;
			ELSE
				CNT_1KHZ <= CNT_1KHZ + 1;
			END IF;
		END IF;
	END PROCESS;
END BEHAV;
