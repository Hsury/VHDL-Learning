--正弦信号发生器 2017/05/08
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SINE_WAVE_GENERATOR IS
	PORT (CLK_50MHZ : IN STD_LOGIC;	--50MHz时钟
	      DATA_OUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));	--量化输出信号
END SINE_WAVE_GENERATOR;

ARCHITECTURE BEHAV OF SINE_WAVE_GENERATOR IS
	COMPONENT WAVE_DATA_ROM IS
	PORT (ADDRESS : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
	      CLOCK : IN STD_LOGIC := '1';
	      Q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
	END COMPONENT;
	
	SIGNAL CNT64 : STD_LOGIC_VECTOR (5 DOWNTO 0);
BEGIN
	PROCESS (CLK_50MHZ)	--6位计数器(索引)
	BEGIN
		IF RISING_EDGE (CLK_50MHZ) THEN
			CNT64 <= CNT64 + 1;	--溢出则自动清零
		END IF;
	END PROCESS;
	
	ROM : WAVE_DATA_ROM PORT MAP (ADDRESS => CNT64,
	                              CLOCK => CLK_50MHZ,
	                              Q => DATA_OUT);
END BEHAV;