--数码管显示模块 2017/04/11
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SEG8 IS
	PORT (DATA_IN : IN INTEGER RANGE 0 TO 9;	--字符输入
	      DP_IN : IN STD_LOGIC;	--小数点输入
	      BAR : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));	--数码管段
END SEG8;

ARCHITECTURE BEHAV OF SEG8 IS
BEGIN
	WITH DATA_IN SELECT
	BAR <= (NOT DP_IN) & "1000000" WHEN 0,
	       (NOT DP_IN) & "1111001" WHEN 1,
	       (NOT DP_IN) & "0100100" WHEN 2,
	       (NOT DP_IN) & "0110000" WHEN 3,
	       (NOT DP_IN) & "0011001" WHEN 4,
	       (NOT DP_IN) & "0010010" WHEN 5,
	       (NOT DP_IN) & "0000010" WHEN 6,
	       (NOT DP_IN) & "1111000" WHEN 7,
	       (NOT DP_IN) & "0000000" WHEN 8,
	       (NOT DP_IN) & "0010000" WHEN 9,
	       "11111111" WHEN OTHERS;
END BEHAV;