--音乐演奏模块 2017/05/11
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MUSIC_BUZZER IS
	PORT (CLK_50MHZ : IN STD_LOGIC;	--50MHz时钟
	      BUZZER : OUT STD_LOGIC);	--无源蜂鸣器
END MUSIC_BUZZER;

ARCHITECTURE BEHAV OF MUSIC_BUZZER IS
	COMPONENT MUSIC_DATA_ROM IS	--LPM_ROM模块
		PORT (ADDRESS : IN STD_LOGIC_VECTOR (10 DOWNTO 0);	--地址
		      CLOCK : IN STD_LOGIC := '1';	--输入端锁存信号
		      Q : OUT STD_LOGIC_VECTOR (8 DOWNTO 0));	--数据
	END COMPONENT;
	
	CONSTANT FREQ_BASS_DO : INTEGER := 262;
	CONSTANT FREQ_BASS_RE : INTEGER := 294;
	CONSTANT FREQ_BASS_MI : INTEGER := 330;
	CONSTANT FREQ_BASS_FA : INTEGER := 349;
	CONSTANT FREQ_BASS_SOL : INTEGER := 392;
	CONSTANT FREQ_BASS_LA : INTEGER := 440;
	CONSTANT FREQ_BASS_TI : INTEGER := 494;
	CONSTANT FREQ_ALTO_DO : INTEGER := 523;
	CONSTANT FREQ_ALTO_RE : INTEGER := 587;
	CONSTANT FREQ_ALTO_MI : INTEGER := 659;
	CONSTANT FREQ_ALTO_FA : INTEGER := 698;
	CONSTANT FREQ_ALTO_SOL : INTEGER := 784;
	CONSTANT FREQ_ALTO_LA : INTEGER := 880;
	CONSTANT FREQ_ALTO_TI : INTEGER := 988;
	CONSTANT FREQ_TREBLE_DO : INTEGER := 1046;
	CONSTANT FREQ_TREBLE_RE : INTEGER := 1175;
	CONSTANT FREQ_TREBLE_MI : INTEGER := 1318;
	CONSTANT FREQ_TREBLE_FA : INTEGER := 1397;
	CONSTANT FREQ_TREBLE_SOL : INTEGER := 1568;
	CONSTANT FREQ_TREBLE_LA : INTEGER := 1760;
	CONSTANT FREQ_TREBLE_TI : INTEGER := 1967;
	
	SIGNAL CNT_BASS_DO : INTEGER RANGE 0 TO (5E7 / FREQ_BASS_DO) - 1;
	SIGNAL CNT_BASS_RE : INTEGER RANGE 0 TO (5E7 / FREQ_BASS_RE) - 1;
	SIGNAL CNT_BASS_MI : INTEGER RANGE 0 TO (5E7 / FREQ_BASS_MI) - 1;
	SIGNAL CNT_BASS_FA : INTEGER RANGE 0 TO (5E7 / FREQ_BASS_FA) - 1;
	SIGNAL CNT_BASS_SOL : INTEGER RANGE 0 TO (5E7 / FREQ_BASS_SOL) - 1;
	SIGNAL CNT_BASS_LA : INTEGER RANGE 0 TO (5E7 / FREQ_BASS_LA) - 1;
	SIGNAL CNT_BASS_TI : INTEGER RANGE 0 TO (5E7 / FREQ_BASS_TI) - 1;
	SIGNAL CNT_ALTO_DO : INTEGER RANGE 0 TO (5E7 / FREQ_ALTO_DO) - 1;
	SIGNAL CNT_ALTO_RE : INTEGER RANGE 0 TO (5E7 / FREQ_ALTO_RE) - 1;
	SIGNAL CNT_ALTO_MI : INTEGER RANGE 0 TO (5E7 / FREQ_ALTO_MI) - 1;
	SIGNAL CNT_ALTO_FA : INTEGER RANGE 0 TO (5E7 / FREQ_ALTO_FA) - 1;
	SIGNAL CNT_ALTO_SOL : INTEGER RANGE 0 TO (5E7 / FREQ_ALTO_SOL) - 1;
	SIGNAL CNT_ALTO_LA : INTEGER RANGE 0 TO (5E7 / FREQ_ALTO_LA) - 1;
	SIGNAL CNT_ALTO_TI : INTEGER RANGE 0 TO (5E7 / FREQ_ALTO_TI) - 1;
	SIGNAL CNT_TREBLE_DO : INTEGER RANGE 0 TO (5E7 / FREQ_TREBLE_DO) - 1;
	SIGNAL CNT_TREBLE_RE : INTEGER RANGE 0 TO (5E7 / FREQ_TREBLE_RE) - 1;
	SIGNAL CNT_TREBLE_MI : INTEGER RANGE 0 TO (5E7 / FREQ_TREBLE_MI) - 1;
	SIGNAL CNT_TREBLE_FA : INTEGER RANGE 0 TO (5E7 / FREQ_TREBLE_FA) - 1;
	SIGNAL CNT_TREBLE_SOL : INTEGER RANGE 0 TO (5E7 / FREQ_TREBLE_SOL) - 1;
	SIGNAL CNT_TREBLE_LA : INTEGER RANGE 0 TO (5E7 / FREQ_TREBLE_LA) - 1;
	SIGNAL CNT_TREBLE_TI : INTEGER RANGE 0 TO (5E7 / FREQ_TREBLE_TI) - 1;
	
	SIGNAL OUTPUT_BASS_DO : STD_LOGIC;
	SIGNAL OUTPUT_BASS_RE : STD_LOGIC;
	SIGNAL OUTPUT_BASS_MI : STD_LOGIC;
	SIGNAL OUTPUT_BASS_FA : STD_LOGIC;
	SIGNAL OUTPUT_BASS_SOL : STD_LOGIC;
	SIGNAL OUTPUT_BASS_LA : STD_LOGIC;
	SIGNAL OUTPUT_BASS_TI : STD_LOGIC;
	SIGNAL OUTPUT_ALTO_DO : STD_LOGIC;
	SIGNAL OUTPUT_ALTO_RE : STD_LOGIC;
	SIGNAL OUTPUT_ALTO_MI : STD_LOGIC;
	SIGNAL OUTPUT_ALTO_FA : STD_LOGIC;
	SIGNAL OUTPUT_ALTO_SOL : STD_LOGIC;
	SIGNAL OUTPUT_ALTO_LA : STD_LOGIC;
	SIGNAL OUTPUT_ALTO_TI : STD_LOGIC;
	SIGNAL OUTPUT_TREBLE_DO : STD_LOGIC;
	SIGNAL OUTPUT_TREBLE_RE : STD_LOGIC;
	SIGNAL OUTPUT_TREBLE_MI : STD_LOGIC;
	SIGNAL OUTPUT_TREBLE_FA : STD_LOGIC;
	SIGNAL OUTPUT_TREBLE_SOL : STD_LOGIC;
	SIGNAL OUTPUT_TREBLE_LA : STD_LOGIC;
	SIGNAL OUTPUT_TREBLE_TI : STD_LOGIC;
	
	CONSTANT CNT_128HZ_OFFSET : INTEGER := 0;	--128Hz时钟计数器补偿值
	
	SIGNAL CLK_128HZ : STD_LOGIC;	--128Hz时钟
	SIGNAL CNT_128HZ : INTEGER RANGE 0 TO 5E7 / (128 - CNT_128HZ_OFFSET) - 1;	--128Hz时钟计数器
	SIGNAL CNT_BEAT : STD_LOGIC_VECTOR (9 DOWNTO 0);	--节拍计数器
	SIGNAL ROM_ADDRESS : STD_LOGIC_VECTOR (10 DOWNTO 0);	--ROM地址
	SIGNAL ROM_DATA : STD_LOGIC_VECTOR (8 DOWNTO 0);	--ROM数据
BEGIN
	ROM : MUSIC_DATA_ROM PORT MAP (ADDRESS => ROM_ADDRESS,
	                               CLOCK => CLK_50MHZ,
	                               Q => ROM_DATA);
	
	PROCESS (CLK_50MHZ)
	BEGIN
		IF RISING_EDGE (CLK_50MHZ) THEN
			CNT_128HZ <= CNT_128HZ + 1;	--128Hz分频器
			IF CNT_128HZ = 0 THEN
				CLK_128HZ <= '1';
			ELSIF CNT_128HZ = 5E7 / (128 - CNT_128HZ_OFFSET) / 2 THEN
				CLK_128HZ <= '0';
			ELSIF CNT_128HZ = 5E7 / (128 - CNT_128HZ_OFFSET) - 1 THEN
				CNT_128HZ <= 0;
			END IF;
			
			CNT_BASS_DO <= CNT_BASS_DO + 1;	--低音Do分频器
			IF CNT_BASS_DO = 0 THEN
				OUTPUT_BASS_DO <= '1';
			ELSIF CNT_BASS_DO = (5E7 / FREQ_BASS_DO) / 2 THEN
				OUTPUT_BASS_DO <= '0';
			ELSIF CNT_BASS_DO = (5E7 / FREQ_BASS_DO) - 1 THEN
				CNT_BASS_DO <= 0;
			END IF;
			
			CNT_BASS_RE <= CNT_BASS_RE + 1;	--低音Re分频器
			IF CNT_BASS_RE = 0 THEN
				OUTPUT_BASS_RE <= '1';
			ELSIF CNT_BASS_RE = (5E7 / FREQ_BASS_RE) / 2 THEN
				OUTPUT_BASS_RE <= '0';
			ELSIF CNT_BASS_RE = (5E7 / FREQ_BASS_RE) - 1 THEN
				CNT_BASS_RE <= 0;
			END IF;
			
			CNT_BASS_MI <= CNT_BASS_MI + 1;	--低音Mi分频器
			IF CNT_BASS_MI = 0 THEN
				OUTPUT_BASS_MI <= '1';
			ELSIF CNT_BASS_MI = (5E7 / FREQ_BASS_MI) / 2 THEN
				OUTPUT_BASS_MI <= '0';
			ELSIF CNT_BASS_MI = (5E7 / FREQ_BASS_MI) - 1 THEN
				CNT_BASS_MI <= 0;
			END IF;
			
			CNT_BASS_FA <= CNT_BASS_FA + 1;	--低音Fa分频器
			IF CNT_BASS_FA = 0 THEN
				OUTPUT_BASS_FA <= '1';
			ELSIF CNT_BASS_FA = (5E7 / FREQ_BASS_FA) / 2 THEN
				OUTPUT_BASS_FA <= '0';
			ELSIF CNT_BASS_FA = (5E7 / FREQ_BASS_FA) - 1 THEN
				CNT_BASS_FA <= 0;
			END IF;
			
			CNT_BASS_SOL <= CNT_BASS_SOL + 1;	--低音Sol分频器
			IF CNT_BASS_SOL = 0 THEN
				OUTPUT_BASS_SOL <= '1';
			ELSIF CNT_BASS_SOL = (5E7 / FREQ_BASS_SOL) / 2 THEN
				OUTPUT_BASS_SOL <= '0';
			ELSIF CNT_BASS_SOL = (5E7 / FREQ_BASS_SOL) - 1 THEN
				CNT_BASS_SOL <= 0;
			END IF;
			
			CNT_BASS_LA <= CNT_BASS_LA + 1;	--低音La分频器
			IF CNT_BASS_LA = 0 THEN
				OUTPUT_BASS_LA <= '1';
			ELSIF CNT_BASS_LA = (5E7 / FREQ_BASS_LA) / 2 THEN
				OUTPUT_BASS_LA <= '0';
			ELSIF CNT_BASS_LA = (5E7 / FREQ_BASS_LA) - 1 THEN
				CNT_BASS_LA <= 0;
			END IF;
			
			CNT_BASS_TI <= CNT_BASS_TI + 1;	--低音Ti分频器
			IF CNT_BASS_TI = 0 THEN
				OUTPUT_BASS_TI <= '1';
			ELSIF CNT_BASS_TI = (5E7 / FREQ_BASS_TI) / 2 THEN
				OUTPUT_BASS_TI <= '0';
			ELSIF CNT_BASS_TI = (5E7 / FREQ_BASS_TI) - 1 THEN
				CNT_BASS_TI <= 0;
			END IF;
			
			CNT_ALTO_DO <= CNT_ALTO_DO + 1;	--中音Do分频器
			IF CNT_ALTO_DO = 0 THEN
				OUTPUT_ALTO_DO <= '1';
			ELSIF CNT_ALTO_DO = (5E7 / FREQ_ALTO_DO) / 2 THEN
				OUTPUT_ALTO_DO <= '0';
			ELSIF CNT_ALTO_DO = (5E7 / FREQ_ALTO_DO) - 1 THEN
				CNT_ALTO_DO <= 0;
			END IF;
			
			CNT_ALTO_RE <= CNT_ALTO_RE + 1;	--中音Re分频器
			IF CNT_ALTO_RE = 0 THEN
				OUTPUT_ALTO_RE <= '1';
			ELSIF CNT_ALTO_RE = (5E7 / FREQ_ALTO_RE) / 2 THEN
				OUTPUT_ALTO_RE <= '0';
			ELSIF CNT_ALTO_RE = (5E7 / FREQ_ALTO_RE) - 1 THEN
				CNT_ALTO_RE <= 0;
			END IF;
			
			CNT_ALTO_MI <= CNT_ALTO_MI + 1;	--中音Mi分频器
			IF CNT_ALTO_MI = 0 THEN
				OUTPUT_ALTO_MI <= '1';
			ELSIF CNT_ALTO_MI = (5E7 / FREQ_ALTO_MI) / 2 THEN
				OUTPUT_ALTO_MI <= '0';
			ELSIF CNT_ALTO_MI = (5E7 / FREQ_ALTO_MI) - 1 THEN
				CNT_ALTO_MI <= 0;
			END IF;
			
			CNT_ALTO_FA <= CNT_ALTO_FA + 1;	--中音Fa分频器
			IF CNT_ALTO_FA = 0 THEN
				OUTPUT_ALTO_FA <= '1';
			ELSIF CNT_ALTO_FA = (5E7 / FREQ_ALTO_FA) / 2 THEN
				OUTPUT_ALTO_FA <= '0';
			ELSIF CNT_ALTO_FA = (5E7 / FREQ_ALTO_FA) - 1 THEN
				CNT_ALTO_FA <= 0;
			END IF;
			
			CNT_ALTO_SOL <= CNT_ALTO_SOL + 1;	--中音Sol分频器
			IF CNT_ALTO_SOL = 0 THEN
				OUTPUT_ALTO_SOL <= '1';
			ELSIF CNT_ALTO_SOL = (5E7 / FREQ_ALTO_SOL) / 2 THEN
				OUTPUT_ALTO_SOL <= '0';
			ELSIF CNT_ALTO_SOL = (5E7 / FREQ_ALTO_SOL) - 1 THEN
				CNT_ALTO_SOL <= 0;
			END IF;
			
			CNT_ALTO_LA <= CNT_ALTO_LA + 1;	--中音La分频器
			IF CNT_ALTO_LA = 0 THEN
				OUTPUT_ALTO_LA <= '1';
			ELSIF CNT_ALTO_LA = (5E7 / FREQ_ALTO_LA) / 2 THEN
				OUTPUT_ALTO_LA <= '0';
			ELSIF CNT_ALTO_LA = (5E7 / FREQ_ALTO_LA) - 1 THEN
				CNT_ALTO_LA <= 0;
			END IF;
			
			CNT_ALTO_TI <= CNT_ALTO_TI + 1;	--中音Ti分频器
			IF CNT_ALTO_TI = 0 THEN
				OUTPUT_ALTO_TI <= '1';
			ELSIF CNT_ALTO_TI = (5E7 / FREQ_ALTO_TI) / 2 THEN
				OUTPUT_ALTO_TI <= '0';
			ELSIF CNT_ALTO_TI = (5E7 / FREQ_ALTO_TI) - 1 THEN
				CNT_ALTO_TI <= 0;
			END IF;
			
			CNT_TREBLE_DO <= CNT_TREBLE_DO + 1;	--高音Do分频器
			IF CNT_TREBLE_DO = 0 THEN
				OUTPUT_TREBLE_DO <= '1';
			ELSIF CNT_TREBLE_DO = (5E7 / FREQ_TREBLE_DO) / 2 THEN
				OUTPUT_TREBLE_DO <= '0';
			ELSIF CNT_TREBLE_DO = (5E7 / FREQ_TREBLE_DO) - 1 THEN
				CNT_TREBLE_DO <= 0;
			END IF;
			
			CNT_TREBLE_RE <= CNT_TREBLE_RE + 1;	--高音Re分频器
			IF CNT_TREBLE_RE = 0 THEN
				OUTPUT_TREBLE_RE <= '1';
			ELSIF CNT_TREBLE_RE = (5E7 / FREQ_TREBLE_RE) / 2 THEN
				OUTPUT_TREBLE_RE <= '0';
			ELSIF CNT_TREBLE_RE = (5E7 / FREQ_TREBLE_RE) - 1 THEN
				CNT_TREBLE_RE <= 0;
			END IF;
			
			CNT_TREBLE_MI <= CNT_TREBLE_MI + 1;	--高音Mi分频器
			IF CNT_TREBLE_MI = 0 THEN
				OUTPUT_TREBLE_MI <= '1';
			ELSIF CNT_TREBLE_MI = (5E7 / FREQ_TREBLE_MI) / 2 THEN
				OUTPUT_TREBLE_MI <= '0';
			ELSIF CNT_TREBLE_MI = (5E7 / FREQ_TREBLE_MI) - 1 THEN
				CNT_TREBLE_MI <= 0;
			END IF;
			
			CNT_TREBLE_FA <= CNT_TREBLE_FA + 1;	--高音Fa分频器
			IF CNT_TREBLE_FA = 0 THEN
				OUTPUT_TREBLE_FA <= '1';
			ELSIF CNT_TREBLE_FA = (5E7 / FREQ_TREBLE_FA) / 2 THEN
				OUTPUT_TREBLE_FA <= '0';
			ELSIF CNT_TREBLE_FA = (5E7 / FREQ_TREBLE_FA) - 1 THEN
				CNT_TREBLE_FA <= 0;
			END IF;
			
			CNT_TREBLE_SOL <= CNT_TREBLE_SOL + 1;	--高音Sol分频器
			IF CNT_TREBLE_SOL = 0 THEN
				OUTPUT_TREBLE_SOL <= '1';
			ELSIF CNT_TREBLE_SOL = (5E7 / FREQ_TREBLE_SOL) / 2 THEN
				OUTPUT_TREBLE_SOL <= '0';
			ELSIF CNT_TREBLE_SOL = (5E7 / FREQ_TREBLE_SOL) - 1 THEN
				CNT_TREBLE_SOL <= 0;
			END IF;
			
			CNT_TREBLE_LA <= CNT_TREBLE_LA + 1;	--高音La分频器
			IF CNT_TREBLE_LA = 0 THEN
				OUTPUT_TREBLE_LA <= '1';
			ELSIF CNT_TREBLE_LA = (5E7 / FREQ_TREBLE_LA) / 2 THEN
				OUTPUT_TREBLE_LA <= '0';
			ELSIF CNT_TREBLE_LA = (5E7 / FREQ_TREBLE_LA) - 1 THEN
				CNT_TREBLE_LA <= 0;
			END IF;
			
			CNT_TREBLE_TI <= CNT_TREBLE_TI + 1;	--高音Ti分频器
			IF CNT_TREBLE_TI = 0 THEN
				OUTPUT_TREBLE_TI <= '1';
			ELSIF CNT_TREBLE_TI = (5E7 / FREQ_TREBLE_TI) / 2 THEN
				OUTPUT_TREBLE_TI <= '0';
			ELSIF CNT_TREBLE_TI = (5E7 / FREQ_TREBLE_TI) - 1 THEN
				CNT_TREBLE_TI <= 0;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (CLK_128HZ)
	BEGIN
		IF RISING_EDGE (CLK_128HZ) THEN
			IF (ROM_DATA = "000000000") THEN	--起始符
				ROM_ADDRESS <= ROM_ADDRESS + 1;
				CNT_BEAT <= (OTHERS => '0');
			ELSIF (ROM_DATA = "111111111") THEN	--终止符
				ROM_ADDRESS <= (OTHERS => '0');
				CNT_BEAT <= (OTHERS => '0');
			ELSE
				IF (ROM_DATA (0) = '0' AND CNT_BEAT = TO_STDLOGICVECTOR ("0000000100" SLL CONV_INTEGER (ROM_DATA (3 DOWNTO 1)))) THEN	--音符断开
					ROM_ADDRESS <= ROM_ADDRESS + 1;
					CNT_BEAT <= (OTHERS => '0');
				ELSIF (ROM_DATA (0) = '1' AND CNT_BEAT = TO_STDLOGICVECTOR ("0000000100" SLL CONV_INTEGER (ROM_DATA (3 DOWNTO 1))) - 1) THEN	--音符连续
					ROM_ADDRESS <= ROM_ADDRESS + 1;
					CNT_BEAT <= (OTHERS => '0');
				ELSE
					CNT_BEAT <= CNT_BEAT + 1;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (ROM_DATA, CNT_BEAT)
	BEGIN
		IF (ROM_DATA (0) = '0' AND CNT_BEAT = TO_STDLOGICVECTOR ("0000000100" SLL CONV_INTEGER (ROM_DATA (3 DOWNTO 1))) - 1) THEN	--添加间隔
			BUZZER <= '0';
		ELSE
			CASE CONV_INTEGER (ROM_DATA (8 DOWNTO 4)) IS
				WHEN 1 => BUZZER <= OUTPUT_BASS_DO;
				WHEN 2 => BUZZER <= OUTPUT_BASS_RE;
				WHEN 3 => BUZZER <= OUTPUT_BASS_MI;
				WHEN 4 => BUZZER <= OUTPUT_BASS_FA;
				WHEN 5 => BUZZER <= OUTPUT_BASS_SOL;
				WHEN 6 => BUZZER <= OUTPUT_BASS_LA;
				WHEN 7 => BUZZER <= OUTPUT_BASS_TI;
				WHEN 8 => BUZZER <= OUTPUT_ALTO_DO;
				WHEN 9 => BUZZER <= OUTPUT_ALTO_RE;
				WHEN 10 => BUZZER <= OUTPUT_ALTO_MI;
				WHEN 11 => BUZZER <= OUTPUT_ALTO_FA;
				WHEN 12 => BUZZER <= OUTPUT_ALTO_SOL;
				WHEN 13 => BUZZER <= OUTPUT_ALTO_LA;
				WHEN 14 => BUZZER <= OUTPUT_ALTO_TI;
				WHEN 15 => BUZZER <= OUTPUT_TREBLE_DO;
				WHEN 16 => BUZZER <= OUTPUT_TREBLE_RE;
				WHEN 17 => BUZZER <= OUTPUT_TREBLE_MI;
				WHEN 18 => BUZZER <= OUTPUT_TREBLE_FA;
				WHEN 19 => BUZZER <= OUTPUT_TREBLE_SOL;
				WHEN 20 => BUZZER <= OUTPUT_TREBLE_LA;
				WHEN 21 => BUZZER <= OUTPUT_TREBLE_TI;
				WHEN OTHERS => BUZZER <= '0';
			END CASE;
		END IF;
	END PROCESS;
END BEHAV;
